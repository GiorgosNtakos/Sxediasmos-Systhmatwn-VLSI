LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
ENTITY testbench4GATES IS
END testbench4GATES;

ARCHITECTURE testbench OF testbench4GATES IS 
    COMPONENT xor8
    GENERIC(
	N: NATURAL :=8);
	PORT(
	 A : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
	 B : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
	 Y : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
	);
	END COMPONENT;
	
	COMPONENT or16
	GENERIC(
	N: NATURAL :=16);
	PORT(
	 A : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
	 B : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
	 Y : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
	);
	END COMPONENT;
	
	COMPONENT nand32
	GENERIC(
	N: NATURAL :=32);
	PORT(
	 A : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
	 B : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
	 Y : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
	);
	END COMPONENT;
	
	COMPONENT nor64
	GENERIC(
	N: NATURAL :=64);
	PORT(
	 A : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
	 B : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
	 Y : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
	);
	END COMPONENT;

	CONSTANT K : NATURAL := 8 ;
	CONSTANT L : NATURAL := 16 ;
	CONSTANT M : NATURAL := 32 ;
	CONSTANT N : NATURAL := 64 ;

	signal ATxor : STD_LOGIC_VECTOR(K-1 DOWNTO 0);
	signal BTxor : STD_LOGIC_VECTOR(K-1 DOWNTO 0);
	signal ATor : STD_LOGIC_VECTOR(L-1 DOWNTO 0);
	signal BTor : STD_LOGIC_VECTOR(L-1 DOWNTO 0);
	signal ATnand : STD_LOGIC_VECTOR(M-1 DOWNTO 0);
	signal BTnand : STD_LOGIC_VECTOR(M-1 DOWNTO 0);
	signal ATnor : STD_LOGIC_VECTOR(N-1 DOWNTO 0);
	signal BTnor : STD_LOGIC_VECTOR(N-1 DOWNTO 0);

	signal YTxor : STD_LOGIC_VECTOR(K-1 DOWNTO 0);
	signal YTor : STD_LOGIC_VECTOR(L-1 DOWNTO 0);
	signal YTnand : STD_LOGIC_VECTOR(M-1 DOWNTO 0);
	signal YTnor : STD_LOGIC_VECTOR(N-1 DOWNTO 0);
	
BEGIN
	
	
	NOR_GATE: nor64 GENERIC MAP(N) PORT MAP(ATnor,BTnor,YTnor);
	NAND_GATE: nand32 GENERIC MAP(M) PORT MAP(ATnand,BTnand,YTnand);
	OR_GATE: or16 GENERIC MAP(L) PORT MAP (ATor,BTor,YTor);
	XOR_GATE: xor8 GENERIC MAP(K) PORT MAP(ATxor,BTxor,YTxor);
	
	stim_proc: process
	BEGIN
	
	ATxor<=X"00";
	BTxor<=X"00";

	ATor<=X"0000";
	BTor<=X"0000";

	ATnand<=X"00000000";
	BTnand<=X"00000000";

	ATnor<=X"0000000000000000";
	BTnor<=X"0000000000000000";
		
		WAIT FOR 20 ns;

	ATxor<=X"00";
	BTxor<=X"FF";

	ATor<=X"0000";
	BTor<=X"FFFF";

	ATnand<=X"00000000";
	BTnand<=X"FFFFFFFF";
		
	ATnor<=X"0000000000000000";
	BTnor<=X"FFFFFFFFFFFFFFFF";
	
		WAIT FOR 20 ns;

	ATxor<=X"FF";
	BTxor<=X"00";

	ATor<=X"FFFF";
	BTor<=X"0000";

	ATnand<=X"FFFFFFFF";
	BTnand<=X"00000000";
		
	ATnor<=X"FFFFFFFFFFFFFFFF";
	BTnor<=X"0000000000000000";
	
		WAIT FOR 20 NS;

	ATxor<=X"FF";
	BTxor<=X"FF";

	ATor<=X"FFFF";
	BTor<=X"FFFF";

	ATnand<=X"FFFFFFFF";
	BTnand<=X"FFFFFFFF";
		
	ATnor<=X"FFFFFFFFFFFFFFFF";
	BTnor<=X"FFFFFFFFFFFFFFFF";
		
		WAIT;
	
	END PROCESS;
	
END;
		
	