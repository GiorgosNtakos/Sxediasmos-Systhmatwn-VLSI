LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

PACKAGE mult_3x3_pack IS

TYPE matrix_in IS ARRAY(NATURAL RANGE <> , NATURAL RANGE <>) OF STD_LOGIC_VECTOR(4 DOWNTO 0);

TYPE matrix_out IS ARRAY(NATURAL RANGE <> , NATURAL RANGE <>) OF STD_LOGIC_VECTOR(9 DOWNTO 0); 

END mult_3x3_pack;