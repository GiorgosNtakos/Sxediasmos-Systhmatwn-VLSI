
LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY bigLunit IS
GENERIC(N: NATURAL :=120);
PORT(

 inp1 : IN std_logic_vector(N-1 DOWNTO 0);
 
 inp2 : IN std_logic_vector(N-1 DOWNTO 0);

 sel  : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
 
 output : OUT std_logic_vector(N-1 DOWNTO 0));
 END bigLunit;
 
 ARCHITECTURE structural OF bigLunit IS
 
 COMPONENT xor8 IS
	GENERIC(N: NATURAL := 8);
	PORT( A : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		  B : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		  Y : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
		  END COMPONENT;
		  
 COMPONENT or16 IS
	GENERIC(N: NATURAL := 16);
	PORT( A : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		  B : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		  Y : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
		  END COMPONENT;
		  
 COMPONENT nand32 IS
	GENERIC(N: NATURAL := 32);
	PORT( A : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		  B : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		  Y : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
		  END COMPONENT;
		  
 COMPONENT nor64 IS
	GENERIC(N: NATURAL := 64);
	PORT( A : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		  B : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		  Y : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
		  END COMPONENT;
		  
COMPONENT mux IS
	GENERIC(N: NATURAL := 8);
	PORT(     a : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		  b : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		  c : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		  d : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		  sel : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		  x : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
		  END COMPONENT;
		  
		  SIGNAL outXor : STD_LOGIC_VECTOR(N-113 DOWNTO 0);
		  SIGNAL outOr : STD_LOGIC_VECTOR(N-97 DOWNTO 8);
		  SIGNAL outNand : STD_LOGIC_VECTOR(N-65 DOWNTO 24);
		  SIGNAL outNOr : STD_LOGIC_VECTOR(N-1 DOWNTO 56);
		  
		  SIGNAl in0_mux : STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		  SIGNAL in1_mux : STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		  SIGNAL in2_mux : STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		  SIGNAL in3_mux : STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		  
BEGIN
 XOR_GATE:  xor8   GENERIC MAP(N-112)  PORT MAP(inp1(N-113 DOWNTO 0),inp2(N-113 DOWNTO 0),outXor);
 OR_GATE:   or16   GENERIC MAP(N-104)  PORT MAP(inp1(N-97 DOWNTO 8),inp2(N-97 DOWNTO 8),outOr);
 NAND_GATE: nand32 GENERIC MAP(N-88)   PORT MAP(inp1(N-65 DOWNTO 24),inp2(N-65 DOWNTO 24),outNand);
 NOR_GATE:  nor64  GENERIC MAP(N-56)   PORT MAP(inp1(N-1 DOWNTO 56),inp2(N-1 DOWNTO 56 ),outNOr);
 
	in0_mux <= (N-1 DOWNTO 8 =>'Z') & outXor;
	in1_mux <= (N-1 DOWNTO 24 =>'Z') & outOr & (7 DOWNTO 0 => 'Z');
	in2_mux <= (N-1 DOWNTO 56 =>'Z') & outNand & (23 DOWNTO 0 =>'Z');
	in3_mux <= outNOr & (55 DOWNTO 0 =>'Z');
 
 
 MUX_GATE: mux     GENERIC MAP(N)      PORT MAP(in0_mux,in1_mux,in2_mux,in3_mux,sel,output);
END structural;